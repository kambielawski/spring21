
package my_package is

	function n_bits_of (X : in integer) return integer;

end package my_package;
